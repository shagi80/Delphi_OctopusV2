�0006586=3000
�0012752=400