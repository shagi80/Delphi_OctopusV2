�0006648=1
�0011945=1
�0006700=1
�0004765=1
�0004766=1
�0005970=1
�0019438=1
�0022371=1
�0006707=1
�0004764=1
�0005971=1